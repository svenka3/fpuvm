// FP-UVM - UVM for FPGAs app 
// Automatically generated from VHDL Package: t_pkg 
package sv_t_pkg; 
  parameter ADDR_W = 16;
  parameter DATA_W = 32;
endpackage : sv_t_pkg 

import sv_t_pkg::* 

